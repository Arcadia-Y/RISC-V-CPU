// Memory Controller
module MemoryController(

);

endmodule