// Data Cache
module DCache(

)

endmodule