// Instruction Cache
module ICache(

)

endmodule