// Reorder Buffer
module ReorderBuffer(

);

endmodule