// Instruction Unit & PC
module InstructionUnit(

);

endmodule