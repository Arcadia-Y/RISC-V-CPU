// Reservation Station & ALU
module ReservationStation(

);

endmodule