// Load Store Buffer
module LoadStoreBuffer(

);

endmodule