// general-purposed cache
module Cache(

)

endmodule