// Register File & Registers
module RegisterFile(

)

endmodule