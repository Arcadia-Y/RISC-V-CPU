// Branch Predictor
module BranchPredictor(

)

endmodule